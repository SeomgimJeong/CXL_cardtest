library ieee;
use ieee.std_logic_1164.all;
package pkg_timestamp is
  -- Constants
  constant TIMESTAMP : std_logic_vector(31 downto 0) := x"69662060";
end pkg_timestamp;
package body pkg_timestamp is
end pkg_timestamp;
